-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"d8080b0b",
    10 => x"0bb5dc08",
    11 => x"0b0b0bb5",
    12 => x"e0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5e00c0b",
    16 => x"0b0bb5dc",
    17 => x"0c0b0b0b",
    18 => x"b5d80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baeec",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5d87080",
    57 => x"c088278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"51889804",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb5e80c",
    65 => x"9f0bb5ec",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b5ec08ff",
    69 => x"05b5ec0c",
    70 => x"b5ec0880",
    71 => x"25eb38b5",
    72 => x"e808ff05",
    73 => x"b5e80cb5",
    74 => x"e8088025",
    75 => x"d738800b",
    76 => x"b5ec0c80",
    77 => x"0bb5e80c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb5e808",
    97 => x"258f3882",
    98 => x"bd2db5e8",
    99 => x"08ff05b5",
   100 => x"e80c82ff",
   101 => x"04b5e808",
   102 => x"b5ec0853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b5e808a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b5ec",
   111 => x"088105b5",
   112 => x"ec0cb5ec",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb5ec0c",
   116 => x"b5e80881",
   117 => x"05b5e80c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b5",
   122 => x"ec088105",
   123 => x"b5ec0cb5",
   124 => x"ec08a02e",
   125 => x"0981068e",
   126 => x"38800bb5",
   127 => x"ec0cb5e8",
   128 => x"088105b5",
   129 => x"e80c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb5f0",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb5f00c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b5",
   169 => x"f0088407",
   170 => x"b5f00c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb290",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b5f00852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b5d80c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d04880b",
   217 => x"ec0c86b7",
   218 => x"2d0402dc",
   219 => x"050d8059",
   220 => x"86e22d81",
   221 => x"0bec0c7a",
   222 => x"52b5f451",
   223 => x"a6a92db5",
   224 => x"d808792e",
   225 => x"80ee38b5",
   226 => x"f80870f8",
   227 => x"0c79ff12",
   228 => x"56595573",
   229 => x"792e8b38",
   230 => x"81187481",
   231 => x"2a555873",
   232 => x"f738f718",
   233 => x"58815980",
   234 => x"752580c8",
   235 => x"38775273",
   236 => x"51848b2d",
   237 => x"b6c052b5",
   238 => x"f451a8df",
   239 => x"2db5d808",
   240 => x"802e9a38",
   241 => x"b6c05783",
   242 => x"fc567670",
   243 => x"84055808",
   244 => x"e80cfc16",
   245 => x"56758025",
   246 => x"f13887e4",
   247 => x"04b5d808",
   248 => x"59848055",
   249 => x"b5f451a8",
   250 => x"b22dfc80",
   251 => x"15811555",
   252 => x"5587a704",
   253 => x"840bec0c",
   254 => x"78802e8d",
   255 => x"38b29451",
   256 => x"8fb72d8d",
   257 => x"ba2d888f",
   258 => x"04b3a851",
   259 => x"8fb72d78",
   260 => x"b5d80c02",
   261 => x"a4050d04",
   262 => x"02f0050d",
   263 => x"840bec0c",
   264 => x"8d882d89",
   265 => x"d72d81f8",
   266 => x"2d83528c",
   267 => x"ed2d8151",
   268 => x"84f02dff",
   269 => x"12527180",
   270 => x"25f13884",
   271 => x"0bec0cb0",
   272 => x"c45185fe",
   273 => x"2d9dc62d",
   274 => x"b5d80880",
   275 => x"2e80f338",
   276 => x"86ea51ae",
   277 => x"e62db294",
   278 => x"518fb72d",
   279 => x"8da72d89",
   280 => x"e32d8fc7",
   281 => x"2db2c00b",
   282 => x"80f52db4",
   283 => x"94087081",
   284 => x"06545553",
   285 => x"71802e85",
   286 => x"38728407",
   287 => x"5373812a",
   288 => x"70810651",
   289 => x"5271802e",
   290 => x"85387288",
   291 => x"07537382",
   292 => x"2a708106",
   293 => x"51527180",
   294 => x"2e853872",
   295 => x"90075373",
   296 => x"832a7081",
   297 => x"06515271",
   298 => x"802e8538",
   299 => x"72a00753",
   300 => x"72fc0c86",
   301 => x"52b5d808",
   302 => x"83388452",
   303 => x"71ec0c88",
   304 => x"df04800b",
   305 => x"b5d80c02",
   306 => x"90050d04",
   307 => x"71980c04",
   308 => x"ffb008b5",
   309 => x"d80c0481",
   310 => x"0bffb00c",
   311 => x"04800bff",
   312 => x"b00c0402",
   313 => x"f4050d8a",
   314 => x"e504b5d8",
   315 => x"0881f02e",
   316 => x"09810689",
   317 => x"38810bb4",
   318 => x"8c0c8ae5",
   319 => x"04b5d808",
   320 => x"81e02e09",
   321 => x"81068938",
   322 => x"810bb490",
   323 => x"0c8ae504",
   324 => x"b5d80852",
   325 => x"b4900880",
   326 => x"2e8838b5",
   327 => x"d8088180",
   328 => x"05527184",
   329 => x"2c728f06",
   330 => x"5353b48c",
   331 => x"08802e99",
   332 => x"38728429",
   333 => x"b3cc0572",
   334 => x"1381712b",
   335 => x"70097308",
   336 => x"06730c51",
   337 => x"53538adb",
   338 => x"04728429",
   339 => x"b3cc0572",
   340 => x"1383712b",
   341 => x"72080772",
   342 => x"0c535380",
   343 => x"0bb4900c",
   344 => x"800bb48c",
   345 => x"0cb68051",
   346 => x"8be62db5",
   347 => x"d808ff24",
   348 => x"fef83880",
   349 => x"0bb5d80c",
   350 => x"028c050d",
   351 => x"0402f805",
   352 => x"0db3cc52",
   353 => x"8f518072",
   354 => x"70840554",
   355 => x"0cff1151",
   356 => x"708025f2",
   357 => x"38028805",
   358 => x"0d0402f0",
   359 => x"050d7551",
   360 => x"89dd2d70",
   361 => x"822cfc06",
   362 => x"b3cc1172",
   363 => x"109e0671",
   364 => x"0870722a",
   365 => x"70830682",
   366 => x"742b7009",
   367 => x"7406760c",
   368 => x"54515657",
   369 => x"53515389",
   370 => x"d72d71b5",
   371 => x"d80c0290",
   372 => x"050d0402",
   373 => x"fc050d72",
   374 => x"5180710c",
   375 => x"800b8412",
   376 => x"0c028405",
   377 => x"0d0402f0",
   378 => x"050d7570",
   379 => x"08841208",
   380 => x"535353ff",
   381 => x"5471712e",
   382 => x"a83889dd",
   383 => x"2d841308",
   384 => x"70842914",
   385 => x"88117008",
   386 => x"7081ff06",
   387 => x"84180881",
   388 => x"11870684",
   389 => x"1a0c5351",
   390 => x"55515151",
   391 => x"89d72d71",
   392 => x"5473b5d8",
   393 => x"0c029005",
   394 => x"0d0402f8",
   395 => x"050d89dd",
   396 => x"2de00870",
   397 => x"8b2a7081",
   398 => x"06515252",
   399 => x"70802e9d",
   400 => x"38b68008",
   401 => x"708429b6",
   402 => x"88057381",
   403 => x"ff06710c",
   404 => x"5151b680",
   405 => x"08811187",
   406 => x"06b6800c",
   407 => x"51800bb6",
   408 => x"a80c89d0",
   409 => x"2d89d72d",
   410 => x"0288050d",
   411 => x"0402fc05",
   412 => x"0d89dd2d",
   413 => x"810bb6a8",
   414 => x"0c89d72d",
   415 => x"b6a80851",
   416 => x"70fa3802",
   417 => x"84050d04",
   418 => x"02fc050d",
   419 => x"b680518b",
   420 => x"d32d8afd",
   421 => x"2d8caa51",
   422 => x"89cc2d02",
   423 => x"84050d04",
   424 => x"b6ac08b5",
   425 => x"d80c0402",
   426 => x"fc050d81",
   427 => x"0bb4980c",
   428 => x"815184f0",
   429 => x"2d028405",
   430 => x"0d0402fc",
   431 => x"050d8dc4",
   432 => x"0489e32d",
   433 => x"80f6518b",
   434 => x"9a2db5d8",
   435 => x"08f33880",
   436 => x"da518b9a",
   437 => x"2db5d808",
   438 => x"e838b5d8",
   439 => x"08b4980c",
   440 => x"b5d80851",
   441 => x"84f02d02",
   442 => x"84050d04",
   443 => x"02ec050d",
   444 => x"76548052",
   445 => x"870b8815",
   446 => x"80f52d56",
   447 => x"53747224",
   448 => x"8338a053",
   449 => x"725182f9",
   450 => x"2d81128b",
   451 => x"1580f52d",
   452 => x"54527272",
   453 => x"25de3802",
   454 => x"94050d04",
   455 => x"02f0050d",
   456 => x"b6ac0854",
   457 => x"81f82d80",
   458 => x"0bb6b00c",
   459 => x"7308802e",
   460 => x"81803882",
   461 => x"0bb5ec0c",
   462 => x"b6b0088f",
   463 => x"06b5e80c",
   464 => x"73085271",
   465 => x"832e9638",
   466 => x"71832689",
   467 => x"3871812e",
   468 => x"af388f9d",
   469 => x"0471852e",
   470 => x"9f388f9d",
   471 => x"04881480",
   472 => x"f52d8415",
   473 => x"08b0dc53",
   474 => x"545285fe",
   475 => x"2d718429",
   476 => x"13700852",
   477 => x"528fa104",
   478 => x"73518dec",
   479 => x"2d8f9d04",
   480 => x"b4940888",
   481 => x"15082c70",
   482 => x"81065152",
   483 => x"71802e87",
   484 => x"38b0e051",
   485 => x"8f9a04b0",
   486 => x"e45185fe",
   487 => x"2d841408",
   488 => x"5185fe2d",
   489 => x"b6b00881",
   490 => x"05b6b00c",
   491 => x"8c14548e",
   492 => x"ac040290",
   493 => x"050d0471",
   494 => x"b6ac0c8e",
   495 => x"9c2db6b0",
   496 => x"08ff05b6",
   497 => x"b40c0402",
   498 => x"e8050db6",
   499 => x"ac08b6b8",
   500 => x"08575580",
   501 => x"f6518b9a",
   502 => x"2db5d808",
   503 => x"812a7081",
   504 => x"06515271",
   505 => x"802ea138",
   506 => x"8fee0489",
   507 => x"e32d80f6",
   508 => x"518b9a2d",
   509 => x"b5d808f3",
   510 => x"38b49808",
   511 => x"813270b4",
   512 => x"980c7052",
   513 => x"5284f02d",
   514 => x"b4980890",
   515 => x"3881fd51",
   516 => x"8b9a2d81",
   517 => x"fa518b9a",
   518 => x"2d95cd04",
   519 => x"81f5518b",
   520 => x"9a2db5d8",
   521 => x"08812a70",
   522 => x"81065152",
   523 => x"71802eaf",
   524 => x"38b6b408",
   525 => x"5271802e",
   526 => x"8938ff12",
   527 => x"b6b40c90",
   528 => x"df04b6b0",
   529 => x"0810b6b0",
   530 => x"08057084",
   531 => x"29165152",
   532 => x"88120880",
   533 => x"2e8938ff",
   534 => x"51881208",
   535 => x"52712d81",
   536 => x"f2518b9a",
   537 => x"2db5d808",
   538 => x"812a7081",
   539 => x"06515271",
   540 => x"802eb138",
   541 => x"b6b008ff",
   542 => x"11b6b408",
   543 => x"56535373",
   544 => x"72258938",
   545 => x"8114b6b4",
   546 => x"0c91a404",
   547 => x"72101370",
   548 => x"84291651",
   549 => x"52881208",
   550 => x"802e8938",
   551 => x"fe518812",
   552 => x"0852712d",
   553 => x"81fd518b",
   554 => x"9a2db5d8",
   555 => x"08812a70",
   556 => x"81065152",
   557 => x"71802ead",
   558 => x"38b6b408",
   559 => x"802e8938",
   560 => x"800bb6b4",
   561 => x"0c91e504",
   562 => x"b6b00810",
   563 => x"b6b00805",
   564 => x"70842916",
   565 => x"51528812",
   566 => x"08802e89",
   567 => x"38fd5188",
   568 => x"12085271",
   569 => x"2d81fa51",
   570 => x"8b9a2db5",
   571 => x"d808812a",
   572 => x"70810651",
   573 => x"5271802e",
   574 => x"ae38b6b0",
   575 => x"08ff1154",
   576 => x"52b6b408",
   577 => x"73258838",
   578 => x"72b6b40c",
   579 => x"92a70471",
   580 => x"10127084",
   581 => x"29165152",
   582 => x"88120880",
   583 => x"2e8938fc",
   584 => x"51881208",
   585 => x"52712db6",
   586 => x"b4087053",
   587 => x"5473802e",
   588 => x"8a388c15",
   589 => x"ff155555",
   590 => x"92ad0482",
   591 => x"0bb5ec0c",
   592 => x"718f06b5",
   593 => x"e80c81eb",
   594 => x"518b9a2d",
   595 => x"b5d80881",
   596 => x"2a708106",
   597 => x"51527180",
   598 => x"2ead3874",
   599 => x"08852e09",
   600 => x"8106a438",
   601 => x"881580f5",
   602 => x"2dff0552",
   603 => x"71881681",
   604 => x"b72d7198",
   605 => x"2b527180",
   606 => x"25883880",
   607 => x"0b881681",
   608 => x"b72d7451",
   609 => x"8dec2d81",
   610 => x"f4518b9a",
   611 => x"2db5d808",
   612 => x"812a7081",
   613 => x"06515271",
   614 => x"802eb338",
   615 => x"7408852e",
   616 => x"098106aa",
   617 => x"38881580",
   618 => x"f52d8105",
   619 => x"52718816",
   620 => x"81b72d71",
   621 => x"81ff068b",
   622 => x"1680f52d",
   623 => x"54527272",
   624 => x"27873872",
   625 => x"881681b7",
   626 => x"2d74518d",
   627 => x"ec2d80da",
   628 => x"518b9a2d",
   629 => x"b5d80881",
   630 => x"2a708106",
   631 => x"51527180",
   632 => x"2e81a638",
   633 => x"b6ac08b6",
   634 => x"b4085553",
   635 => x"73802e8a",
   636 => x"388c13ff",
   637 => x"15555393",
   638 => x"ec047208",
   639 => x"5271822e",
   640 => x"a6387182",
   641 => x"26893871",
   642 => x"812ea938",
   643 => x"95890471",
   644 => x"832eb138",
   645 => x"71842e09",
   646 => x"810680ed",
   647 => x"38881308",
   648 => x"518fb72d",
   649 => x"958904b6",
   650 => x"b4085188",
   651 => x"13085271",
   652 => x"2d958904",
   653 => x"810b8814",
   654 => x"082bb494",
   655 => x"0832b494",
   656 => x"0c94df04",
   657 => x"881380f5",
   658 => x"2d81058b",
   659 => x"1480f52d",
   660 => x"53547174",
   661 => x"24833880",
   662 => x"54738814",
   663 => x"81b72d8e",
   664 => x"9c2d9589",
   665 => x"04750880",
   666 => x"2ea23875",
   667 => x"08518b9a",
   668 => x"2db5d808",
   669 => x"81065271",
   670 => x"802e8b38",
   671 => x"b6b40851",
   672 => x"84160852",
   673 => x"712d8816",
   674 => x"5675da38",
   675 => x"8054800b",
   676 => x"b5ec0c73",
   677 => x"8f06b5e8",
   678 => x"0ca05273",
   679 => x"b6b4082e",
   680 => x"09810698",
   681 => x"38b6b008",
   682 => x"ff057432",
   683 => x"70098105",
   684 => x"7072079f",
   685 => x"2a917131",
   686 => x"51515353",
   687 => x"715182f9",
   688 => x"2d811454",
   689 => x"8e7425c6",
   690 => x"38b49808",
   691 => x"5271b5d8",
   692 => x"0c029805",
   693 => x"0d0402f4",
   694 => x"050dd452",
   695 => x"81ff720c",
   696 => x"71085381",
   697 => x"ff720c72",
   698 => x"882b83fe",
   699 => x"80067208",
   700 => x"7081ff06",
   701 => x"51525381",
   702 => x"ff720c72",
   703 => x"7107882b",
   704 => x"72087081",
   705 => x"ff065152",
   706 => x"5381ff72",
   707 => x"0c727107",
   708 => x"882b7208",
   709 => x"7081ff06",
   710 => x"7207b5d8",
   711 => x"0c525302",
   712 => x"8c050d04",
   713 => x"02f4050d",
   714 => x"74767181",
   715 => x"ff06d40c",
   716 => x"5353b6bc",
   717 => x"08853871",
   718 => x"892b5271",
   719 => x"982ad40c",
   720 => x"71902a70",
   721 => x"81ff06d4",
   722 => x"0c517188",
   723 => x"2a7081ff",
   724 => x"06d40c51",
   725 => x"7181ff06",
   726 => x"d40c7290",
   727 => x"2a7081ff",
   728 => x"06d40c51",
   729 => x"d4087081",
   730 => x"ff065151",
   731 => x"82b8bf52",
   732 => x"7081ff2e",
   733 => x"09810694",
   734 => x"3881ff0b",
   735 => x"d40cd408",
   736 => x"7081ff06",
   737 => x"ff145451",
   738 => x"5171e538",
   739 => x"70b5d80c",
   740 => x"028c050d",
   741 => x"0402fc05",
   742 => x"0d81c751",
   743 => x"81ff0bd4",
   744 => x"0cff1151",
   745 => x"708025f4",
   746 => x"38028405",
   747 => x"0d0402f4",
   748 => x"050d81ff",
   749 => x"0bd40c93",
   750 => x"53805287",
   751 => x"fc80c151",
   752 => x"96a42db5",
   753 => x"d8088b38",
   754 => x"81ff0bd4",
   755 => x"0c815397",
   756 => x"db049795",
   757 => x"2dff1353",
   758 => x"72df3872",
   759 => x"b5d80c02",
   760 => x"8c050d04",
   761 => x"02ec050d",
   762 => x"810bb6bc",
   763 => x"0c8454d0",
   764 => x"08708f2a",
   765 => x"70810651",
   766 => x"515372f3",
   767 => x"3872d00c",
   768 => x"97952db0",
   769 => x"e85185fe",
   770 => x"2dd00870",
   771 => x"8f2a7081",
   772 => x"06515153",
   773 => x"72f33881",
   774 => x"0bd00cb1",
   775 => x"53805284",
   776 => x"d480c051",
   777 => x"96a42db5",
   778 => x"d808812e",
   779 => x"93387282",
   780 => x"2ebd38ff",
   781 => x"135372e5",
   782 => x"38ff1454",
   783 => x"73ffb038",
   784 => x"97952d83",
   785 => x"aa52849c",
   786 => x"80c85196",
   787 => x"a42db5d8",
   788 => x"08812e09",
   789 => x"81069238",
   790 => x"95d62db5",
   791 => x"d80883ff",
   792 => x"ff065372",
   793 => x"83aa2e9d",
   794 => x"3897ae2d",
   795 => x"998004b0",
   796 => x"f45185fe",
   797 => x"2d80539a",
   798 => x"ce04b18c",
   799 => x"5185fe2d",
   800 => x"80549aa0",
   801 => x"0481ff0b",
   802 => x"d40cb154",
   803 => x"97952d8f",
   804 => x"cf538052",
   805 => x"87fc80f7",
   806 => x"5196a42d",
   807 => x"b5d80855",
   808 => x"b5d80881",
   809 => x"2e098106",
   810 => x"9b3881ff",
   811 => x"0bd40c82",
   812 => x"0a52849c",
   813 => x"80e95196",
   814 => x"a42db5d8",
   815 => x"08802e8d",
   816 => x"3897952d",
   817 => x"ff135372",
   818 => x"c9389a93",
   819 => x"0481ff0b",
   820 => x"d40cb5d8",
   821 => x"085287fc",
   822 => x"80fa5196",
   823 => x"a42db5d8",
   824 => x"08b13881",
   825 => x"ff0bd40c",
   826 => x"d4085381",
   827 => x"ff0bd40c",
   828 => x"81ff0bd4",
   829 => x"0c81ff0b",
   830 => x"d40c81ff",
   831 => x"0bd40c72",
   832 => x"862a7081",
   833 => x"06765651",
   834 => x"53729538",
   835 => x"b5d80854",
   836 => x"9aa00473",
   837 => x"822efee2",
   838 => x"38ff1454",
   839 => x"73feed38",
   840 => x"73b6bc0c",
   841 => x"738b3881",
   842 => x"5287fc80",
   843 => x"d05196a4",
   844 => x"2d81ff0b",
   845 => x"d40cd008",
   846 => x"708f2a70",
   847 => x"81065151",
   848 => x"5372f338",
   849 => x"72d00c81",
   850 => x"ff0bd40c",
   851 => x"815372b5",
   852 => x"d80c0294",
   853 => x"050d0402",
   854 => x"e8050d78",
   855 => x"55805681",
   856 => x"ff0bd40c",
   857 => x"d008708f",
   858 => x"2a708106",
   859 => x"51515372",
   860 => x"f3388281",
   861 => x"0bd00c81",
   862 => x"ff0bd40c",
   863 => x"775287fc",
   864 => x"80d15196",
   865 => x"a42d80db",
   866 => x"c6df54b5",
   867 => x"d808802e",
   868 => x"8a38b1ac",
   869 => x"5185fe2d",
   870 => x"9bee0481",
   871 => x"ff0bd40c",
   872 => x"d4087081",
   873 => x"ff065153",
   874 => x"7281fe2e",
   875 => x"0981069d",
   876 => x"3880ff53",
   877 => x"95d62db5",
   878 => x"d8087570",
   879 => x"8405570c",
   880 => x"ff135372",
   881 => x"8025ed38",
   882 => x"81569bd3",
   883 => x"04ff1454",
   884 => x"73c93881",
   885 => x"ff0bd40c",
   886 => x"81ff0bd4",
   887 => x"0cd00870",
   888 => x"8f2a7081",
   889 => x"06515153",
   890 => x"72f33872",
   891 => x"d00c75b5",
   892 => x"d80c0298",
   893 => x"050d0402",
   894 => x"e8050d77",
   895 => x"797b5855",
   896 => x"55805372",
   897 => x"7625a338",
   898 => x"74708105",
   899 => x"5680f52d",
   900 => x"74708105",
   901 => x"5680f52d",
   902 => x"52527171",
   903 => x"2e863881",
   904 => x"519cac04",
   905 => x"8113539c",
   906 => x"83048051",
   907 => x"70b5d80c",
   908 => x"0298050d",
   909 => x"0402ec05",
   910 => x"0d765574",
   911 => x"802ebb38",
   912 => x"9a1580e0",
   913 => x"2d51a9b5",
   914 => x"2db5d808",
   915 => x"b5d808bc",
   916 => x"f00cb5d8",
   917 => x"085454bc",
   918 => x"cc08802e",
   919 => x"99389415",
   920 => x"80e02d51",
   921 => x"a9b52db5",
   922 => x"d808902b",
   923 => x"83fff00a",
   924 => x"06707507",
   925 => x"515372bc",
   926 => x"f00cbcf0",
   927 => x"08537280",
   928 => x"2e9938bc",
   929 => x"c408fe14",
   930 => x"7129bcd8",
   931 => x"0805bcf4",
   932 => x"0c70842b",
   933 => x"bcd00c54",
   934 => x"9dc104bc",
   935 => x"dc08bcf0",
   936 => x"0cbce008",
   937 => x"bcf40cbc",
   938 => x"cc08802e",
   939 => x"8a38bcc4",
   940 => x"08842b53",
   941 => x"9dbd04bc",
   942 => x"e408842b",
   943 => x"5372bcd0",
   944 => x"0c029405",
   945 => x"0d0402d8",
   946 => x"050d800b",
   947 => x"bccc0c84",
   948 => x"5497e42d",
   949 => x"b5d80880",
   950 => x"2e9538b6",
   951 => x"c0528051",
   952 => x"9ad72db5",
   953 => x"d808802e",
   954 => x"8638fe54",
   955 => x"9df704ff",
   956 => x"14547380",
   957 => x"24db3873",
   958 => x"8c38b1bc",
   959 => x"5185fe2d",
   960 => x"7355a380",
   961 => x"04805681",
   962 => x"0bbcf80c",
   963 => x"8853b1d0",
   964 => x"52b6f651",
   965 => x"9bf72db5",
   966 => x"d808762e",
   967 => x"09810687",
   968 => x"38b5d808",
   969 => x"bcf80c88",
   970 => x"53b1dc52",
   971 => x"b792519b",
   972 => x"f72db5d8",
   973 => x"088738b5",
   974 => x"d808bcf8",
   975 => x"0cbcf808",
   976 => x"802e80f6",
   977 => x"38ba860b",
   978 => x"80f52dba",
   979 => x"870b80f5",
   980 => x"2d71982b",
   981 => x"71902b07",
   982 => x"ba880b80",
   983 => x"f52d7088",
   984 => x"2b7207ba",
   985 => x"890b80f5",
   986 => x"2d7107ba",
   987 => x"be0b80f5",
   988 => x"2dbabf0b",
   989 => x"80f52d71",
   990 => x"882b0753",
   991 => x"5f54525a",
   992 => x"56575573",
   993 => x"81abaa2e",
   994 => x"0981068d",
   995 => x"387551a9",
   996 => x"852db5d8",
   997 => x"08569fa6",
   998 => x"047382d4",
   999 => x"d52e8738",
  1000 => x"b1e8519f",
  1001 => x"e704b6c0",
  1002 => x"5275519a",
  1003 => x"d72db5d8",
  1004 => x"0855b5d8",
  1005 => x"08802e83",
  1006 => x"c7388853",
  1007 => x"b1dc52b7",
  1008 => x"92519bf7",
  1009 => x"2db5d808",
  1010 => x"8938810b",
  1011 => x"bccc0c9f",
  1012 => x"ed048853",
  1013 => x"b1d052b6",
  1014 => x"f6519bf7",
  1015 => x"2db5d808",
  1016 => x"802e8a38",
  1017 => x"b1fc5185",
  1018 => x"fe2da0c7",
  1019 => x"04babe0b",
  1020 => x"80f52d54",
  1021 => x"7380d52e",
  1022 => x"09810680",
  1023 => x"ca38babf",
  1024 => x"0b80f52d",
  1025 => x"547381aa",
  1026 => x"2e098106",
  1027 => x"ba38800b",
  1028 => x"b6c00b80",
  1029 => x"f52d5654",
  1030 => x"7481e92e",
  1031 => x"83388154",
  1032 => x"7481eb2e",
  1033 => x"8c388055",
  1034 => x"73752e09",
  1035 => x"810682d0",
  1036 => x"38b6cb0b",
  1037 => x"80f52d55",
  1038 => x"748d38b6",
  1039 => x"cc0b80f5",
  1040 => x"2d547382",
  1041 => x"2e863880",
  1042 => x"55a38004",
  1043 => x"b6cd0b80",
  1044 => x"f52d70bc",
  1045 => x"c40cff05",
  1046 => x"bcc80cb6",
  1047 => x"ce0b80f5",
  1048 => x"2db6cf0b",
  1049 => x"80f52d58",
  1050 => x"76057782",
  1051 => x"80290570",
  1052 => x"bcd40cb6",
  1053 => x"d00b80f5",
  1054 => x"2d70bce8",
  1055 => x"0cbccc08",
  1056 => x"59575876",
  1057 => x"802e81a3",
  1058 => x"388853b1",
  1059 => x"dc52b792",
  1060 => x"519bf72d",
  1061 => x"b5d80881",
  1062 => x"e738bcc4",
  1063 => x"0870842b",
  1064 => x"bcd00c70",
  1065 => x"bce40cb6",
  1066 => x"e50b80f5",
  1067 => x"2db6e40b",
  1068 => x"80f52d71",
  1069 => x"82802905",
  1070 => x"b6e60b80",
  1071 => x"f52d7084",
  1072 => x"80802912",
  1073 => x"b6e70b80",
  1074 => x"f52d7081",
  1075 => x"800a2912",
  1076 => x"70bcec0c",
  1077 => x"bce80871",
  1078 => x"29bcd408",
  1079 => x"0570bcd8",
  1080 => x"0cb6ed0b",
  1081 => x"80f52db6",
  1082 => x"ec0b80f5",
  1083 => x"2d718280",
  1084 => x"2905b6ee",
  1085 => x"0b80f52d",
  1086 => x"70848080",
  1087 => x"2912b6ef",
  1088 => x"0b80f52d",
  1089 => x"70982b81",
  1090 => x"f00a0672",
  1091 => x"0570bcdc",
  1092 => x"0cfe117e",
  1093 => x"297705bc",
  1094 => x"e00c5259",
  1095 => x"5243545e",
  1096 => x"51525952",
  1097 => x"5d575957",
  1098 => x"a2f904b6",
  1099 => x"d20b80f5",
  1100 => x"2db6d10b",
  1101 => x"80f52d71",
  1102 => x"82802905",
  1103 => x"70bcd00c",
  1104 => x"70a02983",
  1105 => x"ff057089",
  1106 => x"2a70bce4",
  1107 => x"0cb6d70b",
  1108 => x"80f52db6",
  1109 => x"d60b80f5",
  1110 => x"2d718280",
  1111 => x"290570bc",
  1112 => x"ec0c7b71",
  1113 => x"291e70bc",
  1114 => x"e00c7dbc",
  1115 => x"dc0c7305",
  1116 => x"bcd80c55",
  1117 => x"5e515155",
  1118 => x"5580519c",
  1119 => x"b52d8155",
  1120 => x"74b5d80c",
  1121 => x"02a8050d",
  1122 => x"0402ec05",
  1123 => x"0d767087",
  1124 => x"2c7180ff",
  1125 => x"06555654",
  1126 => x"bccc088a",
  1127 => x"3873882c",
  1128 => x"7481ff06",
  1129 => x"5455b6c0",
  1130 => x"52bcd408",
  1131 => x"15519ad7",
  1132 => x"2db5d808",
  1133 => x"54b5d808",
  1134 => x"802eb338",
  1135 => x"bccc0880",
  1136 => x"2e983872",
  1137 => x"8429b6c0",
  1138 => x"05700852",
  1139 => x"53a9852d",
  1140 => x"b5d808f0",
  1141 => x"0a0653a3",
  1142 => x"ec047210",
  1143 => x"b6c00570",
  1144 => x"80e02d52",
  1145 => x"53a9b52d",
  1146 => x"b5d80853",
  1147 => x"725473b5",
  1148 => x"d80c0294",
  1149 => x"050d0402",
  1150 => x"e0050d79",
  1151 => x"70842cbc",
  1152 => x"f4080571",
  1153 => x"8f065255",
  1154 => x"53728938",
  1155 => x"b6c05273",
  1156 => x"519ad72d",
  1157 => x"72a029b6",
  1158 => x"c0055480",
  1159 => x"7480f52d",
  1160 => x"56537473",
  1161 => x"2e833881",
  1162 => x"537481e5",
  1163 => x"2e81ef38",
  1164 => x"81707406",
  1165 => x"54587280",
  1166 => x"2e81e338",
  1167 => x"8b1480f5",
  1168 => x"2d70832a",
  1169 => x"79065856",
  1170 => x"769838b4",
  1171 => x"9c085372",
  1172 => x"883872ba",
  1173 => x"c00b81b7",
  1174 => x"2d76b49c",
  1175 => x"0c7353a6",
  1176 => x"a004758f",
  1177 => x"2e098106",
  1178 => x"81b43874",
  1179 => x"9f068d29",
  1180 => x"bab31151",
  1181 => x"53811480",
  1182 => x"f52d7370",
  1183 => x"81055581",
  1184 => x"b72d8314",
  1185 => x"80f52d73",
  1186 => x"70810555",
  1187 => x"81b72d85",
  1188 => x"1480f52d",
  1189 => x"73708105",
  1190 => x"5581b72d",
  1191 => x"871480f5",
  1192 => x"2d737081",
  1193 => x"055581b7",
  1194 => x"2d891480",
  1195 => x"f52d7370",
  1196 => x"81055581",
  1197 => x"b72d8e14",
  1198 => x"80f52d73",
  1199 => x"70810555",
  1200 => x"81b72d90",
  1201 => x"1480f52d",
  1202 => x"73708105",
  1203 => x"5581b72d",
  1204 => x"921480f5",
  1205 => x"2d737081",
  1206 => x"055581b7",
  1207 => x"2d941480",
  1208 => x"f52d7370",
  1209 => x"81055581",
  1210 => x"b72d9614",
  1211 => x"80f52d73",
  1212 => x"70810555",
  1213 => x"81b72d98",
  1214 => x"1480f52d",
  1215 => x"73708105",
  1216 => x"5581b72d",
  1217 => x"9c1480f5",
  1218 => x"2d737081",
  1219 => x"055581b7",
  1220 => x"2d9e1480",
  1221 => x"f52d7381",
  1222 => x"b72d77b4",
  1223 => x"9c0c8053",
  1224 => x"72b5d80c",
  1225 => x"02a0050d",
  1226 => x"0402cc05",
  1227 => x"0d7e605e",
  1228 => x"5a800bbc",
  1229 => x"f008bcf4",
  1230 => x"08595c56",
  1231 => x"8058bcd0",
  1232 => x"08782e81",
  1233 => x"ae38778f",
  1234 => x"06a01757",
  1235 => x"54738f38",
  1236 => x"b6c05276",
  1237 => x"51811757",
  1238 => x"9ad72db6",
  1239 => x"c0568076",
  1240 => x"80f52d56",
  1241 => x"5474742e",
  1242 => x"83388154",
  1243 => x"7481e52e",
  1244 => x"80f63881",
  1245 => x"70750655",
  1246 => x"5c73802e",
  1247 => x"80ea388b",
  1248 => x"1680f52d",
  1249 => x"98065978",
  1250 => x"80de388b",
  1251 => x"537c5275",
  1252 => x"519bf72d",
  1253 => x"b5d80880",
  1254 => x"cf389c16",
  1255 => x"0851a985",
  1256 => x"2db5d808",
  1257 => x"841b0c9a",
  1258 => x"1680e02d",
  1259 => x"51a9b52d",
  1260 => x"b5d808b5",
  1261 => x"d808881c",
  1262 => x"0cb5d808",
  1263 => x"5555bccc",
  1264 => x"08802e98",
  1265 => x"38941680",
  1266 => x"e02d51a9",
  1267 => x"b52db5d8",
  1268 => x"08902b83",
  1269 => x"fff00a06",
  1270 => x"70165154",
  1271 => x"73881b0c",
  1272 => x"787a0c7b",
  1273 => x"54a8a904",
  1274 => x"811858bc",
  1275 => x"d0087826",
  1276 => x"fed438bc",
  1277 => x"cc08802e",
  1278 => x"ae387a51",
  1279 => x"a3892db5",
  1280 => x"d808b5d8",
  1281 => x"0880ffff",
  1282 => x"fff80655",
  1283 => x"5b7380ff",
  1284 => x"fffff82e",
  1285 => x"9238b5d8",
  1286 => x"08fe05bc",
  1287 => x"c40829bc",
  1288 => x"d8080557",
  1289 => x"a6bc0480",
  1290 => x"5473b5d8",
  1291 => x"0c02b405",
  1292 => x"0d0402f4",
  1293 => x"050d7470",
  1294 => x"08810571",
  1295 => x"0c7008bc",
  1296 => x"c8080653",
  1297 => x"53718e38",
  1298 => x"88130851",
  1299 => x"a3892db5",
  1300 => x"d8088814",
  1301 => x"0c810bb5",
  1302 => x"d80c028c",
  1303 => x"050d0402",
  1304 => x"f0050d75",
  1305 => x"881108fe",
  1306 => x"05bcc408",
  1307 => x"29bcd808",
  1308 => x"117208bc",
  1309 => x"c8080605",
  1310 => x"79555354",
  1311 => x"549ad72d",
  1312 => x"0290050d",
  1313 => x"0402f405",
  1314 => x"0d747088",
  1315 => x"2a83fe80",
  1316 => x"06707298",
  1317 => x"2a077288",
  1318 => x"2b87fc80",
  1319 => x"80067398",
  1320 => x"2b81f00a",
  1321 => x"06717307",
  1322 => x"07b5d80c",
  1323 => x"56515351",
  1324 => x"028c050d",
  1325 => x"0402f805",
  1326 => x"0d028e05",
  1327 => x"80f52d74",
  1328 => x"882b0770",
  1329 => x"83ffff06",
  1330 => x"b5d80c51",
  1331 => x"0288050d",
  1332 => x"0402f405",
  1333 => x"0d747678",
  1334 => x"53545280",
  1335 => x"71259738",
  1336 => x"72708105",
  1337 => x"5480f52d",
  1338 => x"72708105",
  1339 => x"5481b72d",
  1340 => x"ff115170",
  1341 => x"eb388072",
  1342 => x"81b72d02",
  1343 => x"8c050d04",
  1344 => x"02e8050d",
  1345 => x"77568070",
  1346 => x"56547376",
  1347 => x"24b138bc",
  1348 => x"d008742e",
  1349 => x"aa387351",
  1350 => x"a3f72db5",
  1351 => x"d808b5d8",
  1352 => x"08098105",
  1353 => x"70b5d808",
  1354 => x"079f2a77",
  1355 => x"05811757",
  1356 => x"57535374",
  1357 => x"76248838",
  1358 => x"bcd00874",
  1359 => x"26d83872",
  1360 => x"b5d80c02",
  1361 => x"98050d04",
  1362 => x"02f0050d",
  1363 => x"b5d40816",
  1364 => x"51aa802d",
  1365 => x"b5d80880",
  1366 => x"2e9b388b",
  1367 => x"53b5d808",
  1368 => x"52bac051",
  1369 => x"a9d12dbc",
  1370 => x"fc085473",
  1371 => x"802e8638",
  1372 => x"bac05173",
  1373 => x"2d029005",
  1374 => x"0d0402dc",
  1375 => x"050d8070",
  1376 => x"5a5574b5",
  1377 => x"d40825af",
  1378 => x"38bcd008",
  1379 => x"752ea838",
  1380 => x"7851a3f7",
  1381 => x"2db5d808",
  1382 => x"09810570",
  1383 => x"b5d80807",
  1384 => x"9f2a7605",
  1385 => x"811b5b56",
  1386 => x"5474b5d4",
  1387 => x"08258838",
  1388 => x"bcd00879",
  1389 => x"26da3880",
  1390 => x"5578bcd0",
  1391 => x"082781cd",
  1392 => x"387851a3",
  1393 => x"f72db5d8",
  1394 => x"08802e81",
  1395 => x"a238b5d8",
  1396 => x"088b0580",
  1397 => x"f52d7084",
  1398 => x"2a708106",
  1399 => x"77107884",
  1400 => x"2bbac00b",
  1401 => x"80f52d5c",
  1402 => x"5c535155",
  1403 => x"5673802e",
  1404 => x"80c63874",
  1405 => x"16822bad",
  1406 => x"b00bb4a8",
  1407 => x"120c5477",
  1408 => x"753110bd",
  1409 => x"80115556",
  1410 => x"90747081",
  1411 => x"055681b7",
  1412 => x"2da07481",
  1413 => x"b72d7681",
  1414 => x"ff068116",
  1415 => x"58547380",
  1416 => x"2e89389c",
  1417 => x"53bac052",
  1418 => x"acb1048b",
  1419 => x"53b5d808",
  1420 => x"52bd8216",
  1421 => x"51ace704",
  1422 => x"7416822b",
  1423 => x"aac80bb4",
  1424 => x"a8120c54",
  1425 => x"7681ff06",
  1426 => x"81165854",
  1427 => x"73802e89",
  1428 => x"389c53ba",
  1429 => x"c052acdf",
  1430 => x"048b53b5",
  1431 => x"d8085277",
  1432 => x"753110bd",
  1433 => x"80055176",
  1434 => x"55a9d12d",
  1435 => x"ad820474",
  1436 => x"90297531",
  1437 => x"7010bd80",
  1438 => x"055154b5",
  1439 => x"d8087481",
  1440 => x"b72d8119",
  1441 => x"59748b24",
  1442 => x"a238abb9",
  1443 => x"04749029",
  1444 => x"75317010",
  1445 => x"bd80058c",
  1446 => x"77315751",
  1447 => x"54807481",
  1448 => x"b72d9e14",
  1449 => x"ff165654",
  1450 => x"74f33802",
  1451 => x"a4050d04",
  1452 => x"02fc050d",
  1453 => x"b5d40813",
  1454 => x"51aa802d",
  1455 => x"b5d80880",
  1456 => x"2e8838b5",
  1457 => x"d808519c",
  1458 => x"b52d800b",
  1459 => x"b5d40caa",
  1460 => x"fa2d8e9c",
  1461 => x"2d028405",
  1462 => x"0d0402fc",
  1463 => x"050d7251",
  1464 => x"70fd2ead",
  1465 => x"3870fd24",
  1466 => x"8a3870fc",
  1467 => x"2e80c438",
  1468 => x"aebb0470",
  1469 => x"fe2eb138",
  1470 => x"70ff2e09",
  1471 => x"8106bc38",
  1472 => x"b5d40851",
  1473 => x"70802eb3",
  1474 => x"38ff11b5",
  1475 => x"d40caebb",
  1476 => x"04b5d408",
  1477 => x"f00570b5",
  1478 => x"d40c5170",
  1479 => x"80259c38",
  1480 => x"800bb5d4",
  1481 => x"0caebb04",
  1482 => x"b5d40881",
  1483 => x"05b5d40c",
  1484 => x"aebb04b5",
  1485 => x"d4089005",
  1486 => x"b5d40caa",
  1487 => x"fa2d8e9c",
  1488 => x"2d028405",
  1489 => x"0d0402fc",
  1490 => x"050d800b",
  1491 => x"b5d40caa",
  1492 => x"fa2d8da0",
  1493 => x"2db5d808",
  1494 => x"b5c40cb4",
  1495 => x"a0518fb7",
  1496 => x"2d028405",
  1497 => x"0d0471bc",
  1498 => x"fc0c0400",
  1499 => x"00ffffff",
  1500 => x"ff00ffff",
  1501 => x"ffff00ff",
  1502 => x"ffffff00",
  1503 => x"4e657074",
  1504 => x"554e4f20",
  1505 => x"534e4553",
  1506 => x"2076302e",
  1507 => x"32000000",
  1508 => x"20202020",
  1509 => x"20202020",
  1510 => x"20202020",
  1511 => x"20202000",
  1512 => x"52657365",
  1513 => x"74000000",
  1514 => x"5363616e",
  1515 => x"6c696e65",
  1516 => x"73000000",
  1517 => x"4a6f7973",
  1518 => x"7469636b",
  1519 => x"20737761",
  1520 => x"70000000",
  1521 => x"50414c00",
  1522 => x"426c656e",
  1523 => x"64000000",
  1524 => x"4c6f6164",
  1525 => x"20524f4d",
  1526 => x"20100000",
  1527 => x"45786974",
  1528 => x"00000000",
  1529 => x"4c6f524f",
  1530 => x"4d206361",
  1531 => x"7274206d",
  1532 => x"61707065",
  1533 => x"72000000",
  1534 => x"4869524f",
  1535 => x"4d206361",
  1536 => x"7274206d",
  1537 => x"61707065",
  1538 => x"72000000",
  1539 => x"45784869",
  1540 => x"526f6d20",
  1541 => x"63617274",
  1542 => x"206d6170",
  1543 => x"70657200",
  1544 => x"4e6f7420",
  1545 => x"73757070",
  1546 => x"6f727465",
  1547 => x"64000000",
  1548 => x"524f4d20",
  1549 => x"6c6f6164",
  1550 => x"20666169",
  1551 => x"6c656400",
  1552 => x"4f4b0000",
  1553 => x"496e6974",
  1554 => x"69616c69",
  1555 => x"7a696e67",
  1556 => x"20534420",
  1557 => x"63617264",
  1558 => x"0a000000",
  1559 => x"16200000",
  1560 => x"14200000",
  1561 => x"15200000",
  1562 => x"53442069",
  1563 => x"6e69742e",
  1564 => x"2e2e0a00",
  1565 => x"53442063",
  1566 => x"61726420",
  1567 => x"72657365",
  1568 => x"74206661",
  1569 => x"696c6564",
  1570 => x"210a0000",
  1571 => x"53444843",
  1572 => x"20657272",
  1573 => x"6f72210a",
  1574 => x"00000000",
  1575 => x"57726974",
  1576 => x"65206661",
  1577 => x"696c6564",
  1578 => x"0a000000",
  1579 => x"52656164",
  1580 => x"20666169",
  1581 => x"6c65640a",
  1582 => x"00000000",
  1583 => x"43617264",
  1584 => x"20696e69",
  1585 => x"74206661",
  1586 => x"696c6564",
  1587 => x"0a000000",
  1588 => x"46415431",
  1589 => x"36202020",
  1590 => x"00000000",
  1591 => x"46415433",
  1592 => x"32202020",
  1593 => x"00000000",
  1594 => x"4e6f2070",
  1595 => x"61727469",
  1596 => x"74696f6e",
  1597 => x"20736967",
  1598 => x"0a000000",
  1599 => x"42616420",
  1600 => x"70617274",
  1601 => x"0a000000",
  1602 => x"4261636b",
  1603 => x"00000000",
  1604 => x"00000002",
  1605 => x"00000002",
  1606 => x"0000177c",
  1607 => x"00000000",
  1608 => x"00000002",
  1609 => x"00001790",
  1610 => x"00000000",
  1611 => x"00000002",
  1612 => x"000017a0",
  1613 => x"0000034e",
  1614 => x"00000003",
  1615 => x"00001998",
  1616 => x"00000004",
  1617 => x"00000001",
  1618 => x"000017a8",
  1619 => x"00000000",
  1620 => x"00000001",
  1621 => x"000017b4",
  1622 => x"00000001",
  1623 => x"00000001",
  1624 => x"000017c4",
  1625 => x"00000002",
  1626 => x"00000001",
  1627 => x"000017c8",
  1628 => x"00000003",
  1629 => x"00000002",
  1630 => x"000017d0",
  1631 => x"00001746",
  1632 => x"00000002",
  1633 => x"000017dc",
  1634 => x"000006ba",
  1635 => x"00000000",
  1636 => x"00000000",
  1637 => x"00000000",
  1638 => x"000017e4",
  1639 => x"000017f8",
  1640 => x"0000180c",
  1641 => x"00001820",
  1642 => x"00000004",
  1643 => x"00001830",
  1644 => x"000019a8",
  1645 => x"00000004",
  1646 => x"00001840",
  1647 => x"00001914",
  1648 => x"00000000",
  1649 => x"00000000",
  1650 => x"00000000",
  1651 => x"00000000",
  1652 => x"00000000",
  1653 => x"00000000",
  1654 => x"00000000",
  1655 => x"00000000",
  1656 => x"00000000",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000002",
  1673 => x"00001e80",
  1674 => x"00001548",
  1675 => x"00000002",
  1676 => x"00001e9e",
  1677 => x"00001548",
  1678 => x"00000002",
  1679 => x"00001ebc",
  1680 => x"00001548",
  1681 => x"00000002",
  1682 => x"00001eda",
  1683 => x"00001548",
  1684 => x"00000002",
  1685 => x"00001ef8",
  1686 => x"00001548",
  1687 => x"00000002",
  1688 => x"00001f16",
  1689 => x"00001548",
  1690 => x"00000002",
  1691 => x"00001f34",
  1692 => x"00001548",
  1693 => x"00000002",
  1694 => x"00001f52",
  1695 => x"00001548",
  1696 => x"00000002",
  1697 => x"00001f70",
  1698 => x"00001548",
  1699 => x"00000002",
  1700 => x"00001f8e",
  1701 => x"00001548",
  1702 => x"00000002",
  1703 => x"00001fac",
  1704 => x"00001548",
  1705 => x"00000002",
  1706 => x"00001fca",
  1707 => x"00001548",
  1708 => x"00000002",
  1709 => x"00001fe8",
  1710 => x"00001548",
  1711 => x"00000004",
  1712 => x"00001908",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
  1716 => x"000016da",
  1717 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

